-- hello_world_qsys.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity hello_world_qsys is
	port (
		button1_external_connection_export : in  std_logic                    := '0'; -- button1_external_connection.export
		button2_external_connection_export : in  std_logic                    := '0'; -- button2_external_connection.export
		button3_external_connection_export : in  std_logic                    := '0'; -- button3_external_connection.export
		button4_external_connection_export : in  std_logic                    := '0'; -- button4_external_connection.export
		clk_clk                            : in  std_logic                    := '0'; --                         clk.clk
		leds_external_connection_export    : out std_logic_vector(4 downto 0);        --    leds_external_connection.export
		reset_reset_n                      : in  std_logic                    := '0'; --                       reset.reset_n
		seg1_external_connection_export    : out std_logic_vector(6 downto 0);        --    seg1_external_connection.export
		seg2_external_connection_export    : out std_logic_vector(6 downto 0);        --    seg2_external_connection.export
		seg3_external_connection_export    : out std_logic_vector(6 downto 0);        --    seg3_external_connection.export
		seg4_external_connection_export    : out std_logic_vector(6 downto 0);        --    seg4_external_connection.export
		seg5_external_connection_export    : out std_logic_vector(6 downto 0);        --    seg5_external_connection.export
		seg6_external_connection_export    : out std_logic_vector(6 downto 0);        --    seg6_external_connection.export
		switch_external_connection_export  : in  std_logic                    := '0'  --  switch_external_connection.export
	);
end entity hello_world_qsys;

architecture rtl of hello_world_qsys is
	component hello_world_qsys_button1 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component hello_world_qsys_button1;

	component hello_world_qsys_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component hello_world_qsys_jtag_uart;

	component hello_world_qsys_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(4 downto 0)                      -- export
		);
	end component hello_world_qsys_leds;

	component hello_world_qsys_nios is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(15 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(15 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component hello_world_qsys_nios;

	component hello_world_qsys_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component hello_world_qsys_ram;

	component hello_world_qsys_seg1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component hello_world_qsys_seg1;

	component hello_world_qsys_mm_interconnect_0 is
		port (
			clk_clk_clk                             : in  std_logic                     := 'X';             -- clk
			nios_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			seg2_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			nios_data_master_address                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			nios_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios_data_master_read                   : in  std_logic                     := 'X';             -- read
			nios_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			nios_data_master_write                  : in  std_logic                     := 'X';             -- write
			nios_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			nios_instruction_master_address         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			nios_instruction_master_read            : in  std_logic                     := 'X';             -- read
			nios_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			button1_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			button1_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button2_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			button2_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button3_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			button3_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button4_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			button4_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			leds_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                           : out std_logic;                                        -- write
			leds_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                      : out std_logic;                                        -- chipselect
			nios_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			nios_debug_mem_slave_write              : out std_logic;                                        -- write
			nios_debug_mem_slave_read               : out std_logic;                                        -- read
			nios_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			nios_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			nios_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			nios_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			ram_s1_address                          : out std_logic_vector(11 downto 0);                    -- address
			ram_s1_write                            : out std_logic;                                        -- write
			ram_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ram_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			ram_s1_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			ram_s1_chipselect                       : out std_logic;                                        -- chipselect
			ram_s1_clken                            : out std_logic;                                        -- clken
			seg1_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			seg1_s1_write                           : out std_logic;                                        -- write
			seg1_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg1_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			seg1_s1_chipselect                      : out std_logic;                                        -- chipselect
			seg2_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			seg2_s1_write                           : out std_logic;                                        -- write
			seg2_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg2_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			seg2_s1_chipselect                      : out std_logic;                                        -- chipselect
			seg3_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			seg3_s1_write                           : out std_logic;                                        -- write
			seg3_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg3_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			seg3_s1_chipselect                      : out std_logic;                                        -- chipselect
			seg4_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			seg4_s1_write                           : out std_logic;                                        -- write
			seg4_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg4_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			seg4_s1_chipselect                      : out std_logic;                                        -- chipselect
			seg5_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			seg5_s1_write                           : out std_logic;                                        -- write
			seg5_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg5_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			seg5_s1_chipselect                      : out std_logic;                                        -- chipselect
			seg6_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			seg6_s1_write                           : out std_logic;                                        -- write
			seg6_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			seg6_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			seg6_s1_chipselect                      : out std_logic;                                        -- chipselect
			switch_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			switch_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component hello_world_qsys_mm_interconnect_0;

	component hello_world_qsys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component hello_world_qsys_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios_debug_reset_request_reset                                : std_logic;                     -- nios:debug_reset_request -> [mm_interconnect_0:seg2_reset_reset_bridge_in_reset_reset, nios_debug_reset_request_reset:in, rst_controller:reset_in1]
	signal nios_data_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	signal nios_data_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	signal nios_data_master_debugaccess                                  : std_logic;                     -- nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	signal nios_data_master_address                                      : std_logic_vector(15 downto 0); -- nios:d_address -> mm_interconnect_0:nios_data_master_address
	signal nios_data_master_byteenable                                   : std_logic_vector(3 downto 0);  -- nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	signal nios_data_master_read                                         : std_logic;                     -- nios:d_read -> mm_interconnect_0:nios_data_master_read
	signal nios_data_master_write                                        : std_logic;                     -- nios:d_write -> mm_interconnect_0:nios_data_master_write
	signal nios_data_master_writedata                                    : std_logic_vector(31 downto 0); -- nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	signal nios_instruction_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	signal nios_instruction_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	signal nios_instruction_master_address                               : std_logic_vector(15 downto 0); -- nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	signal nios_instruction_master_read                                  : std_logic;                     -- nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_nios_debug_mem_slave_readdata               : std_logic_vector(31 downto 0); -- nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	signal mm_interconnect_0_nios_debug_mem_slave_waitrequest            : std_logic;                     -- nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios_debug_mem_slave_debugaccess            : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios_debug_mem_slave_address                : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	signal mm_interconnect_0_nios_debug_mem_slave_read                   : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	signal mm_interconnect_0_nios_debug_mem_slave_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios_debug_mem_slave_write                  : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	signal mm_interconnect_0_nios_debug_mem_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	signal mm_interconnect_0_ram_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	signal mm_interconnect_0_ram_s1_readdata                             : std_logic_vector(31 downto 0); -- ram:readdata -> mm_interconnect_0:ram_s1_readdata
	signal mm_interconnect_0_ram_s1_address                              : std_logic_vector(11 downto 0); -- mm_interconnect_0:ram_s1_address -> ram:address
	signal mm_interconnect_0_ram_s1_byteenable                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	signal mm_interconnect_0_ram_s1_write                                : std_logic;                     -- mm_interconnect_0:ram_s1_write -> ram:write
	signal mm_interconnect_0_ram_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:ram_s1_writedata -> ram:writedata
	signal mm_interconnect_0_ram_s1_clken                                : std_logic;                     -- mm_interconnect_0:ram_s1_clken -> ram:clken
	signal mm_interconnect_0_seg1_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:seg1_s1_chipselect -> seg1:chipselect
	signal mm_interconnect_0_seg1_s1_readdata                            : std_logic_vector(31 downto 0); -- seg1:readdata -> mm_interconnect_0:seg1_s1_readdata
	signal mm_interconnect_0_seg1_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:seg1_s1_address -> seg1:address
	signal mm_interconnect_0_seg1_s1_write                               : std_logic;                     -- mm_interconnect_0:seg1_s1_write -> mm_interconnect_0_seg1_s1_write:in
	signal mm_interconnect_0_seg1_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:seg1_s1_writedata -> seg1:writedata
	signal mm_interconnect_0_seg2_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:seg2_s1_chipselect -> seg2:chipselect
	signal mm_interconnect_0_seg2_s1_readdata                            : std_logic_vector(31 downto 0); -- seg2:readdata -> mm_interconnect_0:seg2_s1_readdata
	signal mm_interconnect_0_seg2_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:seg2_s1_address -> seg2:address
	signal mm_interconnect_0_seg2_s1_write                               : std_logic;                     -- mm_interconnect_0:seg2_s1_write -> mm_interconnect_0_seg2_s1_write:in
	signal mm_interconnect_0_seg2_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:seg2_s1_writedata -> seg2:writedata
	signal mm_interconnect_0_seg3_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:seg3_s1_chipselect -> seg3:chipselect
	signal mm_interconnect_0_seg3_s1_readdata                            : std_logic_vector(31 downto 0); -- seg3:readdata -> mm_interconnect_0:seg3_s1_readdata
	signal mm_interconnect_0_seg3_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:seg3_s1_address -> seg3:address
	signal mm_interconnect_0_seg3_s1_write                               : std_logic;                     -- mm_interconnect_0:seg3_s1_write -> mm_interconnect_0_seg3_s1_write:in
	signal mm_interconnect_0_seg3_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:seg3_s1_writedata -> seg3:writedata
	signal mm_interconnect_0_seg4_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:seg4_s1_chipselect -> seg4:chipselect
	signal mm_interconnect_0_seg4_s1_readdata                            : std_logic_vector(31 downto 0); -- seg4:readdata -> mm_interconnect_0:seg4_s1_readdata
	signal mm_interconnect_0_seg4_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:seg4_s1_address -> seg4:address
	signal mm_interconnect_0_seg4_s1_write                               : std_logic;                     -- mm_interconnect_0:seg4_s1_write -> mm_interconnect_0_seg4_s1_write:in
	signal mm_interconnect_0_seg4_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:seg4_s1_writedata -> seg4:writedata
	signal mm_interconnect_0_seg5_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:seg5_s1_chipselect -> seg5:chipselect
	signal mm_interconnect_0_seg5_s1_readdata                            : std_logic_vector(31 downto 0); -- seg5:readdata -> mm_interconnect_0:seg5_s1_readdata
	signal mm_interconnect_0_seg5_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:seg5_s1_address -> seg5:address
	signal mm_interconnect_0_seg5_s1_write                               : std_logic;                     -- mm_interconnect_0:seg5_s1_write -> mm_interconnect_0_seg5_s1_write:in
	signal mm_interconnect_0_seg5_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:seg5_s1_writedata -> seg5:writedata
	signal mm_interconnect_0_seg6_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:seg6_s1_chipselect -> seg6:chipselect
	signal mm_interconnect_0_seg6_s1_readdata                            : std_logic_vector(31 downto 0); -- seg6:readdata -> mm_interconnect_0:seg6_s1_readdata
	signal mm_interconnect_0_seg6_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:seg6_s1_address -> seg6:address
	signal mm_interconnect_0_seg6_s1_write                               : std_logic;                     -- mm_interconnect_0:seg6_s1_write -> mm_interconnect_0_seg6_s1_write:in
	signal mm_interconnect_0_seg6_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:seg6_s1_writedata -> seg6:writedata
	signal mm_interconnect_0_switch_s1_readdata                          : std_logic_vector(31 downto 0); -- switch:readdata -> mm_interconnect_0:switch_s1_readdata
	signal mm_interconnect_0_switch_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_s1_address -> switch:address
	signal mm_interconnect_0_button1_s1_readdata                         : std_logic_vector(31 downto 0); -- button1:readdata -> mm_interconnect_0:button1_s1_readdata
	signal mm_interconnect_0_button1_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button1_s1_address -> button1:address
	signal mm_interconnect_0_button2_s1_readdata                         : std_logic_vector(31 downto 0); -- button2:readdata -> mm_interconnect_0:button2_s1_readdata
	signal mm_interconnect_0_button2_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button2_s1_address -> button2:address
	signal mm_interconnect_0_button3_s1_readdata                         : std_logic_vector(31 downto 0); -- button3:readdata -> mm_interconnect_0:button3_s1_readdata
	signal mm_interconnect_0_button3_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button3_s1_address -> button3:address
	signal mm_interconnect_0_button4_s1_readdata                         : std_logic_vector(31 downto 0); -- button4:readdata -> mm_interconnect_0:button4_s1_readdata
	signal mm_interconnect_0_button4_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button4_s1_address -> button4:address
	signal mm_interconnect_0_leds_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                            : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                               : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal nios_irq_irq                                                  : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [nios:reset_req, ram:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal nios_debug_reset_request_reset_ports_inv                      : std_logic;                     -- nios_debug_reset_request_reset:inv -> [button1:reset_n, button2:reset_n, button3:reset_n, button4:reset_n, leds:reset_n, seg2:reset_n, seg3:reset_n, seg4:reset_n, seg5:reset_n, seg6:reset_n, switch:reset_n]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_seg1_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_seg1_s1_write:inv -> seg1:write_n
	signal mm_interconnect_0_seg2_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_seg2_s1_write:inv -> seg2:write_n
	signal mm_interconnect_0_seg3_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_seg3_s1_write:inv -> seg3:write_n
	signal mm_interconnect_0_seg4_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_seg4_s1_write:inv -> seg4:write_n
	signal mm_interconnect_0_seg5_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_seg5_s1_write:inv -> seg5:write_n
	signal mm_interconnect_0_seg6_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_seg6_s1_write:inv -> seg6:write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag_uart:rst_n, nios:reset_n, seg1:reset_n]

begin

	button1 : component hello_world_qsys_button1
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => nios_debug_reset_request_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_button1_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_button1_s1_readdata,    --                    .readdata
			in_port  => button1_external_connection_export        -- external_connection.export
		);

	button2 : component hello_world_qsys_button1
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => nios_debug_reset_request_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_button2_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_button2_s1_readdata,    --                    .readdata
			in_port  => button2_external_connection_export        -- external_connection.export
		);

	button3 : component hello_world_qsys_button1
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => nios_debug_reset_request_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_button3_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_button3_s1_readdata,    --                    .readdata
			in_port  => button3_external_connection_export        -- external_connection.export
		);

	button4 : component hello_world_qsys_button1
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => nios_debug_reset_request_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_button4_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_button4_s1_readdata,    --                    .readdata
			in_port  => button4_external_connection_export        -- external_connection.export
		);

	jtag_uart : component hello_world_qsys_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	leds : component hello_world_qsys_leds
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => nios_debug_reset_request_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_external_connection_export            -- external_connection.export
		);

	nios : component hello_world_qsys_nios
		port map (
			clk                                 => clk_clk,                                            --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,           --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                 --                          .reset_req
			d_address                           => nios_data_master_address,                           --               data_master.address
			d_byteenable                        => nios_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios_data_master_read,                              --                          .read
			d_readdata                          => nios_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios_data_master_write,                             --                          .write
			d_writedata                         => nios_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios_instruction_master_read,                       --                          .read
			i_readdata                          => nios_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                -- custom_instruction_master.readra
		);

	ram : component hello_world_qsys_ram
		port map (
			clk        => clk_clk,                             --   clk1.clk
			address    => mm_interconnect_0_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,  --       .reset_req
			freeze     => '0'                                  -- (terminated)
		);

	seg1 : component hello_world_qsys_seg1
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_seg1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seg1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seg1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seg1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seg1_s1_readdata,        --                    .readdata
			out_port   => seg1_external_connection_export            -- external_connection.export
		);

	seg2 : component hello_world_qsys_seg1
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => nios_debug_reset_request_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_seg2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seg2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seg2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seg2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seg2_s1_readdata,        --                    .readdata
			out_port   => seg2_external_connection_export            -- external_connection.export
		);

	seg3 : component hello_world_qsys_seg1
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => nios_debug_reset_request_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_seg3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seg3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seg3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seg3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seg3_s1_readdata,        --                    .readdata
			out_port   => seg3_external_connection_export            -- external_connection.export
		);

	seg4 : component hello_world_qsys_seg1
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => nios_debug_reset_request_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_seg4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seg4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seg4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seg4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seg4_s1_readdata,        --                    .readdata
			out_port   => seg4_external_connection_export            -- external_connection.export
		);

	seg5 : component hello_world_qsys_seg1
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => nios_debug_reset_request_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_seg5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seg5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seg5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seg5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seg5_s1_readdata,        --                    .readdata
			out_port   => seg5_external_connection_export            -- external_connection.export
		);

	seg6 : component hello_world_qsys_seg1
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => nios_debug_reset_request_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_seg6_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_seg6_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_seg6_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_seg6_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_seg6_s1_readdata,        --                    .readdata
			out_port   => seg6_external_connection_export            -- external_connection.export
		);

	switch : component hello_world_qsys_button1
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => nios_debug_reset_request_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_switch_s1_readdata,     --                    .readdata
			in_port  => switch_external_connection_export         -- external_connection.export
		);

	mm_interconnect_0 : component hello_world_qsys_mm_interconnect_0
		port map (
			clk_clk_clk                             => clk_clk,                                                   --                          clk_clk.clk
			nios_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                            -- nios_reset_reset_bridge_in_reset.reset
			seg2_reset_reset_bridge_in_reset_reset  => nios_debug_reset_request_reset,                            -- seg2_reset_reset_bridge_in_reset.reset
			nios_data_master_address                => nios_data_master_address,                                  --                 nios_data_master.address
			nios_data_master_waitrequest            => nios_data_master_waitrequest,                              --                                 .waitrequest
			nios_data_master_byteenable             => nios_data_master_byteenable,                               --                                 .byteenable
			nios_data_master_read                   => nios_data_master_read,                                     --                                 .read
			nios_data_master_readdata               => nios_data_master_readdata,                                 --                                 .readdata
			nios_data_master_write                  => nios_data_master_write,                                    --                                 .write
			nios_data_master_writedata              => nios_data_master_writedata,                                --                                 .writedata
			nios_data_master_debugaccess            => nios_data_master_debugaccess,                              --                                 .debugaccess
			nios_instruction_master_address         => nios_instruction_master_address,                           --          nios_instruction_master.address
			nios_instruction_master_waitrequest     => nios_instruction_master_waitrequest,                       --                                 .waitrequest
			nios_instruction_master_read            => nios_instruction_master_read,                              --                                 .read
			nios_instruction_master_readdata        => nios_instruction_master_readdata,                          --                                 .readdata
			button1_s1_address                      => mm_interconnect_0_button1_s1_address,                      --                       button1_s1.address
			button1_s1_readdata                     => mm_interconnect_0_button1_s1_readdata,                     --                                 .readdata
			button2_s1_address                      => mm_interconnect_0_button2_s1_address,                      --                       button2_s1.address
			button2_s1_readdata                     => mm_interconnect_0_button2_s1_readdata,                     --                                 .readdata
			button3_s1_address                      => mm_interconnect_0_button3_s1_address,                      --                       button3_s1.address
			button3_s1_readdata                     => mm_interconnect_0_button3_s1_readdata,                     --                                 .readdata
			button4_s1_address                      => mm_interconnect_0_button4_s1_address,                      --                       button4_s1.address
			button4_s1_readdata                     => mm_interconnect_0_button4_s1_readdata,                     --                                 .readdata
			jtag_uart_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --      jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                 .write
			jtag_uart_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                 .read
			jtag_uart_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                 .readdata
			jtag_uart_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                 .writedata
			jtag_uart_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                 .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                 .chipselect
			leds_s1_address                         => mm_interconnect_0_leds_s1_address,                         --                          leds_s1.address
			leds_s1_write                           => mm_interconnect_0_leds_s1_write,                           --                                 .write
			leds_s1_readdata                        => mm_interconnect_0_leds_s1_readdata,                        --                                 .readdata
			leds_s1_writedata                       => mm_interconnect_0_leds_s1_writedata,                       --                                 .writedata
			leds_s1_chipselect                      => mm_interconnect_0_leds_s1_chipselect,                      --                                 .chipselect
			nios_debug_mem_slave_address            => mm_interconnect_0_nios_debug_mem_slave_address,            --             nios_debug_mem_slave.address
			nios_debug_mem_slave_write              => mm_interconnect_0_nios_debug_mem_slave_write,              --                                 .write
			nios_debug_mem_slave_read               => mm_interconnect_0_nios_debug_mem_slave_read,               --                                 .read
			nios_debug_mem_slave_readdata           => mm_interconnect_0_nios_debug_mem_slave_readdata,           --                                 .readdata
			nios_debug_mem_slave_writedata          => mm_interconnect_0_nios_debug_mem_slave_writedata,          --                                 .writedata
			nios_debug_mem_slave_byteenable         => mm_interconnect_0_nios_debug_mem_slave_byteenable,         --                                 .byteenable
			nios_debug_mem_slave_waitrequest        => mm_interconnect_0_nios_debug_mem_slave_waitrequest,        --                                 .waitrequest
			nios_debug_mem_slave_debugaccess        => mm_interconnect_0_nios_debug_mem_slave_debugaccess,        --                                 .debugaccess
			ram_s1_address                          => mm_interconnect_0_ram_s1_address,                          --                           ram_s1.address
			ram_s1_write                            => mm_interconnect_0_ram_s1_write,                            --                                 .write
			ram_s1_readdata                         => mm_interconnect_0_ram_s1_readdata,                         --                                 .readdata
			ram_s1_writedata                        => mm_interconnect_0_ram_s1_writedata,                        --                                 .writedata
			ram_s1_byteenable                       => mm_interconnect_0_ram_s1_byteenable,                       --                                 .byteenable
			ram_s1_chipselect                       => mm_interconnect_0_ram_s1_chipselect,                       --                                 .chipselect
			ram_s1_clken                            => mm_interconnect_0_ram_s1_clken,                            --                                 .clken
			seg1_s1_address                         => mm_interconnect_0_seg1_s1_address,                         --                          seg1_s1.address
			seg1_s1_write                           => mm_interconnect_0_seg1_s1_write,                           --                                 .write
			seg1_s1_readdata                        => mm_interconnect_0_seg1_s1_readdata,                        --                                 .readdata
			seg1_s1_writedata                       => mm_interconnect_0_seg1_s1_writedata,                       --                                 .writedata
			seg1_s1_chipselect                      => mm_interconnect_0_seg1_s1_chipselect,                      --                                 .chipselect
			seg2_s1_address                         => mm_interconnect_0_seg2_s1_address,                         --                          seg2_s1.address
			seg2_s1_write                           => mm_interconnect_0_seg2_s1_write,                           --                                 .write
			seg2_s1_readdata                        => mm_interconnect_0_seg2_s1_readdata,                        --                                 .readdata
			seg2_s1_writedata                       => mm_interconnect_0_seg2_s1_writedata,                       --                                 .writedata
			seg2_s1_chipselect                      => mm_interconnect_0_seg2_s1_chipselect,                      --                                 .chipselect
			seg3_s1_address                         => mm_interconnect_0_seg3_s1_address,                         --                          seg3_s1.address
			seg3_s1_write                           => mm_interconnect_0_seg3_s1_write,                           --                                 .write
			seg3_s1_readdata                        => mm_interconnect_0_seg3_s1_readdata,                        --                                 .readdata
			seg3_s1_writedata                       => mm_interconnect_0_seg3_s1_writedata,                       --                                 .writedata
			seg3_s1_chipselect                      => mm_interconnect_0_seg3_s1_chipselect,                      --                                 .chipselect
			seg4_s1_address                         => mm_interconnect_0_seg4_s1_address,                         --                          seg4_s1.address
			seg4_s1_write                           => mm_interconnect_0_seg4_s1_write,                           --                                 .write
			seg4_s1_readdata                        => mm_interconnect_0_seg4_s1_readdata,                        --                                 .readdata
			seg4_s1_writedata                       => mm_interconnect_0_seg4_s1_writedata,                       --                                 .writedata
			seg4_s1_chipselect                      => mm_interconnect_0_seg4_s1_chipselect,                      --                                 .chipselect
			seg5_s1_address                         => mm_interconnect_0_seg5_s1_address,                         --                          seg5_s1.address
			seg5_s1_write                           => mm_interconnect_0_seg5_s1_write,                           --                                 .write
			seg5_s1_readdata                        => mm_interconnect_0_seg5_s1_readdata,                        --                                 .readdata
			seg5_s1_writedata                       => mm_interconnect_0_seg5_s1_writedata,                       --                                 .writedata
			seg5_s1_chipselect                      => mm_interconnect_0_seg5_s1_chipselect,                      --                                 .chipselect
			seg6_s1_address                         => mm_interconnect_0_seg6_s1_address,                         --                          seg6_s1.address
			seg6_s1_write                           => mm_interconnect_0_seg6_s1_write,                           --                                 .write
			seg6_s1_readdata                        => mm_interconnect_0_seg6_s1_readdata,                        --                                 .readdata
			seg6_s1_writedata                       => mm_interconnect_0_seg6_s1_writedata,                       --                                 .writedata
			seg6_s1_chipselect                      => mm_interconnect_0_seg6_s1_chipselect,                      --                                 .chipselect
			switch_s1_address                       => mm_interconnect_0_switch_s1_address,                       --                        switch_s1.address
			switch_s1_readdata                      => mm_interconnect_0_switch_s1_readdata                       --                                 .readdata
		);

	irq_mapper : component hello_world_qsys_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios_irq_irq                    --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => nios_debug_reset_request_reset,     -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	nios_debug_reset_request_reset_ports_inv <= not nios_debug_reset_request_reset;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_seg1_s1_write_ports_inv <= not mm_interconnect_0_seg1_s1_write;

	mm_interconnect_0_seg2_s1_write_ports_inv <= not mm_interconnect_0_seg2_s1_write;

	mm_interconnect_0_seg3_s1_write_ports_inv <= not mm_interconnect_0_seg3_s1_write;

	mm_interconnect_0_seg4_s1_write_ports_inv <= not mm_interconnect_0_seg4_s1_write;

	mm_interconnect_0_seg5_s1_write_ports_inv <= not mm_interconnect_0_seg5_s1_write;

	mm_interconnect_0_seg6_s1_write_ports_inv <= not mm_interconnect_0_seg6_s1_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of hello_world_qsys
